/*
   CS/ECE 552 Spring '22
  
   Filename        : decode.v
   Description     : This is the module for the overall decode stage of the processor.
*/
`default_nettype none
module decode (/* TODO: Add appropriate inputs/outputs for your decode stage here*/);

   wire immSrc;
   wire ALUJump;
   wire MemWrt;
   wire InvA;
   wire InvB;
   wire Cin;
   wire sign;
   wire brType;
   wire BSrc;
   wire 0ext;
   wire ALUOpr;
   wire RegDst;
   wire RegSrc;
   wire RegWrt;

      

endmodule
`default_nettype wire
